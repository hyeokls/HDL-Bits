module top_module (
    input [7:0] a,
    input [7:0] b,
    output [7:0] s,
    output overflow
); 
    
    assign s = a+b;
    assign overflow = (a[7] & b[7] & ~s[7]) | (~a[7] & ~b[7] & s[7] );

endmodule

00000_0010  +2
00111_1111  +127
01000_0001  +129
01111_1110  +254

01111_1111  -127
01000_0001  -1
11000_0000  -128
11111_1110  -254

01000_0001
01000_0001
10000_0010

0_0101_1010
0_0101_1010
0_1011_0100 

